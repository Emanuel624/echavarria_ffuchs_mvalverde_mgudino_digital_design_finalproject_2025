module dmem (
  input  logic        clk,
  input  logic        we,
  input  logic [31:0] a, wd,
  output logic [31:0] rd
);
  // 64 palabras de 32 bits: índices 0..63
  logic [31:0] RAM [0:63];

  // Lectura combinacional (word-aligned).
  // Para 64 palabras usamos 6 bits de índice: a[7:2]
  assign rd = RAM[a[7:2]];

  // Escritura sincrónica
  always_ff @(posedge clk) begin
    if (we) RAM[a[7:2]] <= wd;
  end
endmodule
