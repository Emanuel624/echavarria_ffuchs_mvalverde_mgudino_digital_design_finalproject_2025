
module alu (
  input  logic [31:0] A,
  input  logic [31:0] B,
  input  logic [1:0]  ALUControl,   // 00=ADD, 01=SUB, 10=AND, 11=ORR
  output logic [31:0] Result,
  output logic [3:0]  ALUFlags      // {N,Z,C,V}
);
  // Internos
  logic [31:0] sum_add, sum_sub;
  logic        c_add, c_sub;
  logic        n, z, c, v;

  // ADD (A + B)
  logic [32:0] add33;
  assign add33   = {1'b0, A} + {1'b0, B};
  assign sum_add = add33[31:0];
  assign c_add   = add33[32];  // carry-out

  // SUB (A - B) = A + (~B) + 1
  logic [32:0] sub33;
  assign sub33   = {1'b0, A} + {1'b0, ~B} + 33'd1;
  assign sum_sub = sub33[31:0];
  assign c_sub   = sub33[32];  // en ARM, C = NOT borrow = carry-out de esta suma

  // Resultado según operación
  always_comb begin
    unique case (ALUControl)
      2'b00: Result = sum_add;        // ADD
      2'b01: Result = sum_sub;        // SUB
      2'b10: Result = (A & B);        // AND
      2'b11: Result = (A | B);        // ORR
      default: Result = 32'b0;
    endcase
  end

  // Flags
  // N: bit 31 del resultado
  // Z: resultado == 0
  // C,V: dependen de la operación (para AND/ORR se ponen 0; el reg de flags decide si se escriben vía FlagW)
  always_comb begin
    n = Result[31];
    z = (Result == 32'b0);

    unique case (ALUControl)
      2'b00: begin // ADD
        c = c_add;
        // overflow en suma con signo: mismos signos en A y B, cambia signo en resultado
        v = (A[31] == B[31]) && (Result[31] != A[31]);
      end
      2'b01: begin // SUB
        c = c_sub; // NOT borrow
        // overflow en resta: signos opuestos entre A y B, cambia signo en resultado
        v = (A[31] != B[31]) && (Result[31] != A[31]);
      end
      default: begin // AND / ORR
        c = 1'b0;
        v = 1'b0;
      end
    endcase
  end

  assign ALUFlags = {n, z, c, v};

endmodule
